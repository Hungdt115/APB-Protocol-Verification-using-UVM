ahskjakjskajkskskj:
